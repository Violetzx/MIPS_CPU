module data_forward(
				
				
				);
endmodule